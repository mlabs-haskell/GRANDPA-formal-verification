Require Import Blocks.AnyBlock.
Require Import Votes.
Require Import State.
Require Import Time.
Require Import RoundNumber.
Require Import Preliminars.
Require Import DataTypes.List.Count.
Require Import DataTypes.List.Fold.
Require Import Protocol.FinalizedBlock.
Require Import Protocol.Io.
Require Import Protocol.Protocol.

Require Import PeanoNat.

Require Import Classes.Functor.
Require Import Classes.Eqb.
Require Import Classes.Math.All.
Require Import Instances.List.

Require Protocol.Proofs.Consistency.old_consistency.
Require Protocol.Proofs.Consistency.Rounds.Existence.
Require Protocol.Proofs.Consistency.Finalization.SubmmiterFinalized.

Open Scope bool.
Open Scope list.
Open Scope eqb.
Open Scope math.
Open Scope natWrapper.

Require Import Lia.

Definition VoterVotedInRound (v:Voter) (opaque:OpaqueRound.OpaqueRoundState)
:Prop
  :=
    (Votes.voter_voted_in_votes v (OpaqueRound.get_all_prevote_votes opaque) = true)
    \/
    (Votes.voter_voted_in_votes v (OpaqueRound.get_all_precommit_votes opaque) = true).

Definition voter_is_hones_at_round `{Io} (v:Voter) (r:RoundNumber) : bool
  :=
  (0 <? count v (get_round_honest_voters r))%nat.


(*
  TODO: Add a module to Finalization called [SubmitterIsParticipant]
that proofs that all finalizations are done by a participant of
   the protocol and move this lemma there
*)
Lemma theorem_4_1_eq_aux `{Io}
(t:Time)
  (fb: FinalizedBlock)
  (b1_in:List.In fb (global_finalized_blocks (get_state_up_to t)))
  :
  exists
  (vr:OpaqueRound.OpaqueRoundState)
  (vr2:OpaqueRound.OpaqueRoundState)
  ,
  let v := fb.(FinalizedBlock.submitter_voter)
  in
    (
      State.get_voter_opaque_round
        (get_state_up_to fb.(FinalizedBlock.time) )
        v
        fb.(FinalizedBlock.round_number)
      =
      Some vr
    )
    /\
    (
      g
        (OpaqueRound.get_all_precommit_votes vr)
      =
      Some fb.(FinalizedBlock.block)
    )
  /\
    (
      State.get_voter_opaque_round
        (get_state_up_to (t+(Time.from_nat 2)*global_time_constant))
        v
        fb.(FinalizedBlock.round_number)
      =
      Some vr2
    ).
Proof.
  Admitted.
  (*
  pose (finalized_block_time_leq b1 round_finalized t1 t b1_in) as t1_leq_t.
  remember (t+(Time.from_nat 2)*global_time_constant) as new_t eqn:new_t_eq.
  assert (List.In (to_any b1,t1, round_finalized) (global_finalized_blocks (get_state_up_to new_t))) as b1_in_new_t.
  {
    pose (finalized_blocks_monotone_over_time2 t (new_t - t) (to_any b1, t1,round_finalized) b1_in).
    enough ((new_t - t +t) = new_t) as H0.
    rewrite <- H0.
    assumption.
    admit.
    (* lia. *)
    }
  destruct (finalized_block_came_from_voter b1 round_finalized t1 new_t  b1_in_new_t) as [v [vr [is_some_vr g_vr]]].
  exists v.
  pose (round_continuos_existence v t1 round_finalized vr is_some_vr (new_t - t1)) as vr_exists_at_new_t.
  assert (new_t - t1 +t1 = new_t) as is_new_t. admit. (* lia. *)
  Admitted.
  *)
  (*
  rewrite is_new_t in vr_exists_at_new_t.
  simpl in vr_exists_at_new_t.
  destruct vr_exists_at_new_t as [vr2 is_some_vr2].
  exists vr.
  exists vr2.
  auto.
Qed.
   *)


Lemma theorem_4_1_eq `{io:Io}
  (t:Time)
  (fb1 fb2 : FinalizedBlock)
  (un_related:
    Unrelated
      fb1.(FinalizedBlock.block).(AnyBlock.block)
      fb2.(FinalizedBlock.block).(AnyBlock.block)
  )
  (fb1_in:List.In fb1 (global_finalized_blocks (get_state_up_to t)))
  (fb2_in:List.In fb2 (global_finalized_blocks (get_state_up_to t)))
  (finalized_same_round : fb1.(FinalizedBlock.round_number) = fb2.(FinalizedBlock.round_number))
  :
  exists
    (t3:Time)
    (v:Voter)
    (r:OpaqueRound.OpaqueRoundState)
    (s:Sets.DictionarySet Voter)
    ,
    (
      (
        Rounds.Existence.IsRoundAt v t3 fb1.(FinalizedBlock.round_number) r
      )
      /\
      (
        List.length (Sets.to_list s)
        >=
        1+ Voters.calculate_max_bizantiners (OpaqueRound.get_prevote_voters r)
      )%nat
      /\
      (forall v2, List.In v2 (Sets.to_list s) -> VoterVotedInRound v2 r)
      /\
      (forall v3, List.In v3 (Sets.to_list s) -> List.In v3 (get_round_bizantine_voters fb1.(FinalizedBlock.round_number) ))
    ).
Proof.
  (**
    We are going to prove that the voter who finalized the  block [fb1]
     at t + synchronisation can see block [fb2] as finalized and has enough
     information to find the set of byzantine voters.
    Why t+synchronisation time?
    To have [fb1] and [fb2] as finalized blocks, we
      must have that [t > max(fb1.time,fb2.time) ]
    So, after synchronisation time we guaranteed that the voter who finalized
     [fb1] can see the finalization information of [fb2].
    We can state this in the lemma explicitly, but is easier to apply it
     in the main theorem if leave it as `exists t3` instead.

  *)
  remember (t + (Time.from_nat 2) * global_time_constant) as new_t eqn:new_t_eq.
  exists new_t.
  remember fb1.(FinalizedBlock.submitter_voter) as v.
  remember fb1.(FinalizedBlock.round_number) as r_n.
  exists v.
  (*
  First step, proof that at t + synchronisation time, the voter of [fb1] has
     a [RoundState].
  In the paper this isn't needed, but without this, we can begin the proof.
  *)
  assert (exists r, Rounds.Existence.IsRoundAt v new_t r_n r).
  {
    (*Proof that [fb1.submitter_voter] has a voter state at the
        finalization time [fb1.time]
      TODO: remove this part definign has_vs, not needed anymore
    *)
    pose (SubmmiterFinalized.finalized_block_was_submitted fb1 fb1_in) as was_finalized.
    destruct was_finalized as [ vs_initial [ r_finalization (vs_is_participant & r_is_at_t1 & in_finalization_list)  ] ].
    assert (forall t, exists vs, get_voter_state v (get_state_up_to t) = Some vs) as has_vs.
    {
      eapply VoterStateExists.participants_has_voter_state_always.
      unfold VoterStateExists.IsParticipant.
      exists vs_initial.
      subst v.
      assumption.
    }

    (*Proof that [v] (the voter who submitted fb1) was a participant of round 0
      this is a basic requirement of a lot of Consistency lemmas.
      *)
    assert (VoterStateExists.IsParticipant v) as has_vs_at_init.
    {
      subst v.
      unfold VoterStateExists.IsParticipant.
      eauto.
    }

    (*
      We have a lemma that allow us to conclude the existence of the round that we want.
      TODO: assert first that fb1.time <= t and fb2.time <= 2
    *)
    pose (Rounds.Existence.continuous_existence has_vs_at_init t ((Time.from_nat 2) * global_time_constant) r_n) as e.
    simpl in e.
    rewrite new_t_eq.
    simpl.
    apply e.
    clear e.
    remember (t - fb1.(FinalizedBlock.time) :Time) as t_increment.
    assert ( t = fb1.(FinalizedBlock.time) + t_increment) as H.
    {
      subst t_increment.
      destruct (fb1.(FinalizedBlock.time)) as [nt_fb1] eqn:fb1_t_eq.
      simpl.
      destruct t as [nt_t] eqn:t_eq.
      simpl.
      enough (nt_t = nt_fb1 + (nt_t - nt_fb1))%nat as H .
      rewrite H at 1. auto.
      apply Arith_base.le_plus_minus_stt.
      pose (Finalization.SubmmiterFinalized.in_finalization_list_means_time_is_at_least _ fb1_in) as H.
      rewrite fb1_t_eq in H.
      simpl in H.
      lia.
    }
    rewrite H.
    clear H.
    eapply (Rounds.Existence.continuous_existence has_vs_at_init fb1.(FinalizedBlock.time) t_increment r_n).
    subst v.
    subst r_n.
    eauto.
  }
  destruct H as [r H].
  exists r.
Qed.

  (*
  remember (t + (Time.from_nat 2) * global_time_constant) as new_t eqn:new_t_eq.
  exists new_t.
  destruct (theorem_4_1_eq_aux b1 round_finalized t1 t b1_in) as [v [v1r [v1r2 [is_some_v1r [g_v1r is_some_v1r2]]]]].
  exists v.
  exists v1r2.
  remember (List.filter (fun v3 => Votes.voter_voted_in_votes v3 (OpaqueRound.get_all_precommit_votes v1r2)) (get_round_bizantine_voters round_finalized)) as s_as_list eqn:s_as_list_eq.
  remember (Sets.from_list s_as_list) as s.
  exists s.
  rewrite <- new_t_eq in is_some_v1r2.
  split.
  assumption.
  split.
  - destruct (theorem_4_1_eq_aux b2 round_finalized t2 t b2_in) as [v2 [v2r [v2r2 [is_some_v2r [g_v2r is_some_v2r2]]]]].
  *)
    (*
       TODO in 3.8 :
       we need to show that after t+2*global_time_constant v has got all the votes on v2r, and as such we have
       a supermajority for both blocks in this round (b1 and b2) at this time.
       Then we destruct the Votes.is_safe predicate applied in the precommits at time t + 2*global_time_constant
       In the False case, we end this sub-proof.
       In the True case, b_1 and b_2 are related by a lemma in the Votes.v about supermajority on safe sets, contra with un_related
    *)
  (*
    The other two parts to be proved, are a consequency of the construction of the list (literally they are in the predicate that build the list).
   *)
    Admitted.



Lemma theorem_4_1_lt `{io:Io}
  (t:Time)
  (fb1 fb2 : FinalizedBlock)
  (un_related:
    Unrelated
      fb1.(FinalizedBlock.block).(AnyBlock.block)
      fb2.(FinalizedBlock.block).(AnyBlock.block)
  )
  (fb1_in:List.In fb1 (global_finalized_blocks (get_state_up_to t)))
  (fb2_in:List.In fb2 (global_finalized_blocks (get_state_up_to t)))
  (symmetry_hipotesis:
    fb1.(FinalizedBlock.round_number)
    <
    fb2.(FinalizedBlock.round_number)
  )
  :
  exists
    (t3:Time)
    (v:Voter)
    (r_n:RoundNumber)
    (r:OpaqueRound.OpaqueRoundState)
    (s:Sets.DictionarySet Voter)
    ,
    (
      (
        Rounds.Existence.IsRoundAt v t3 r_n r
      )
      /\
      (
        List.length (Sets.to_list s)
        >=
        1+ Voters.calculate_max_bizantiners (OpaqueRound.get_prevote_voters r)
      )%nat
      /\
      (forall v2, List.In v2 (Sets.to_list s) -> VoterVotedInRound v2 r)
      /\
      (forall v3, List.In v3 (Sets.to_list s) -> List.In v3 (get_round_bizantine_voters r_n))
    ).
Proof.
  (*
  dependent induction b1.
  - pose (originBlock_is_always_prefix b2) as contra.
    apply (prefix_implies_related _ _) in contra.
    contradiction.
  - dependent destruction b2.
    +  pose (originBlock_is_always_prefix (NewBlock b1 id)) as contra.
       apply (prefix_implies_related _ _) in contra.
       apply related_symmetric in contra.
       contradiction.
    +
      (*TODO in 3.8 *)
  *)
Admitted.


(** Theorem 4.1
The original lemma states that

  if we finalized two unrelated blocks
  [fb1] y [fb1], then we can find a set [s] of voters such that
     |s| >= 1
  and all of the voters in [s] voted in a particular vote. Even better
  there exists a synchronous way to find such a set.

This doesn't tell anything a bout a synchronous procedure,
but by virtue of coq constructive logic, the proof
of this theorem shows the existence of a procedure to
find the set.

Additionally, we need to state the theorem conclusion in
terms of the particular view of a particular voter at some time.
This, since we don't have a notion of
  " all the votes emitted for a round at a time"
ad
*)
Theorem theorem_4_1 `{io:Io}
  (t:Time)
  (fb1 fb2 : FinalizedBlock)
  (un_related:
    Unrelated
      fb1.(FinalizedBlock.block).(AnyBlock.block)
      fb2.(FinalizedBlock.block).(AnyBlock.block)
  )
  (fb1_in:
    List.In fb1 (global_finalized_blocks (get_state_up_to t))
  )
  (fb2_in:
    List.In fb2 (global_finalized_blocks (get_state_up_to t))
  )
  :
  exists
    (t3:Time)
    (v:Voter)
    (r_n:RoundNumber)
    (r:OpaqueRound.OpaqueRoundState)
    (s:Sets.DictionarySet Voter)
    ,
    (
      ((* Exists a voter [v] that sees the round [r] at time [t3].
          All the rest of the statements reference to the view of
          this particular voter v.
      *)
        Rounds.Existence.IsRoundAt v t3 r_n r
      )
      /\
      ((* Exists a set [s] with at least [1+f] voters of round [r].*)
        List.length (Sets.to_list s)
        >=
        1+ Voters.calculate_max_bizantiners (OpaqueRound.get_prevote_voters r)
      )%nat
      /\
      (*  All voters of  [s] emitted a vote  in round [r]. *)
      (forall v2, List.In v2 (Sets.to_list s) -> VoterVotedInRound v2 r)
      /\
      (* All voters of [s] are byzantine voters for round [r] *)
      (forall v3, List.In v3 (Sets.to_list s) -> List.In v3 (get_round_bizantine_voters r_n))
    ).
Proof.
  (* Use naturals trichotomy to stablish for [fb1] y [fb2] tree possible cases:
     - fb1 was finalized in a round below fb2
     - fb1 and fb2 where finalized in the same round
     - fb2 was finalized in a round below fb1.
     Name this fact as [trico]
  *)
  pose (
    Arith.Compare_dec.lt_eq_lt_dec
    (RoundNumber.to_nat fb1.(FinalizedBlock.round_number))
    (RoundNumber.to_nat fb2.(FinalizedBlock.round_number))
  ) as trico.
  (* Tell the interpreter we are going to handle the tree cases
     by separate and rename trico according to the hypothesis.
  *)
  destruct trico as [[fb1_n_lt_fb2_n | fb1_n_eq_fb2_n]| fb2_n_lt_fb1_n].
  (*Solve the case fb1 finalized in a round below fb2, by using lemma
     [theorem_4_1_lt] for it.
  *)
  - apply (
      theorem_4_1_lt
        t
        fb1
        fb2
        un_related
        fb1_in
        fb2_in
        fb1_n_lt_fb2_n
    );try assumption.
  (* Focus on case for fb1 and fb2 finalized in the same round.*)
  -
    (* Convince coq that we can apply our auxiliar theorem here*)
    assert( fb1.(round_number) = fb2.(round_number) ) as fb1_n_eq_fb2_n_2. {
      destruct (fb1.(round_number)).
      destruct (fb2.(round_number)).
      auto.
    }
    (* Applying [theorem_4_1_eq] for this case*)
    destruct (
      theorem_4_1_eq
        t
        fb1
        fb2
        un_related
        fb1_in
        fb2_in
        fb1_n_eq_fb2_n_2
    ) as [t3 [v3 [ r [s result]]]].
    exists t3.
    exists v3.
    exists (fb1.(FinalizedBlock.round_number)).
    exists r.
    exists s.
    assumption.
    (*Focus case fb2 was finalized in a round below fb1 *)
  -
    (*Telling coq that the fact that two blocks are unrelated is symmetric*)
    pose (
      Blocks.Block.unrelated_symmetric
        fb1.(block).(AnyBlock.block)
        fb2.(block).(AnyBlock.block)
        un_related
    ) as un_related2.
    (*Solving this case by using theorem_4_1_lt*)
    apply (
      theorem_4_1_lt
      t
      fb2
      fb1
      un_related2
      fb2_in
      fb1_in
    );try assumption.
Qed.


Corollary corollary_4_3
  `{Io}
  (round_finalized_number:RoundNumber)
  (time_finalied:Time)
  (b_finalized:AnyBlock)
  (v:Voter)
  (r_n:RoundNumber)
  (is_honest: voter_is_hones_at_round v r_n = true)
  (t_increment:Time)
  (r_n_geq: r_n >= round_finalized_number)
  (opaque_r_n : OpaqueRound.OpaqueRoundState)
  (opaque_from_state
    :
    State.get_voter_opaque_round (get_state_up_to (t_increment + time_finalied) ) v r_n
    = Some opaque_r_n
  )
  (r_n_completable:
   OpaqueRound.is_completable opaque_r_n = true
  )
  :exists (eb:AnyBlock),
    (
      OpaqueRound.get_estimate opaque_r_n
      =
      Some eb
    )
    /\
    (
      Block.is_prefix b_finalized.(AnyBlock.block) eb.(AnyBlock.block) = true
    ).
Proof.
  (*TODO: delayed until 3.8
   *)
  Admitted.

Close Scope bool.
Close Scope list.
Close Scope eqb.
Close Scope math.
Close Scope natWrapper.
